module register_select();
    
endmodule